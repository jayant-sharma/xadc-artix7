module adc_12bit()

port din;


//test suraj demo
endmodule
